LIBRARY IEEE;
USE IEEE.STD_logic_1164.all;

ENTITY fulladder is
port(
  a: in std_logic;
  b: in std_logic;
  cin: in std_logic;
  s: out std_logic;
  cout: out std_logic
);
end fulladder;

architecture arq_fulladder of fulladder is
begin
  s <= a xor b xor cin;
  cout <= (a and b) or (a and cin) or (b and cin);
end arq_fulladder;