------------------------------------------------------------------------------------------
-- FILENAME:  fpu.vhd
-- TITLE: Floating Point Unit
-- PROJECT: 
-- PURPOSE: Top module
-- VERSION: 
-- AUTHOR: David Cemin
-- DATE:   Sat 26 May 2012 06:03:00 PM BRT
------------------------------------------------------------------------------------------

------------------------------------------------------------------------------------------
--Libraries
------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;


------------------------------------------------------------------------------------------
--Entity
------------------------------------------------------------------------------------------
entity fpu is
	port(
		);
end entity;

------------------------------------------------------------------------------------------
--Architecture
------------------------------------------------------------------------------------------
architecture fpu of fpu is


		------------------------------------------
		-- Types
		------------------------------------------


		------------------------------------------
		-- Constants
		------------------------------------------


		------------------------------------------
		-- Signal Declarations
		------------------------------------------


begin


		------------------------------------------
		-- Port Mappings
		------------------------------------------


		------------------------------------------
		-- Processes
		------------------------------------------


		------------------------------------------
		-- Asynchronous Assignments
		------------------------------------------


end fpu;

