LIBRARY IEEE;
USE  IEEE.STD_LOGIC_1164.all;
USE  IEEE.STD_LOGIC_ARITH.all;
USE  IEEE.STD_LOGIC_UNSIGNED.all;
-- This code displays time in the DE2's LCD Display
-- Key2  resets time
ENTITY Operativa IS
PORT(
  reset, clk, btn0, btn1, btn2: IN STD_LOGIC;
  DATA_BUS: INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
  LCD_RW: BUFFER STD_LOGIC;
  LCD_RS, LCD_E, LCD_ON, RESET_LED: OUT STD_LOGIC;
  
  word_data_in, posicao0, posicao1: in std_logic_vector(3 downto 0);
  reg_data_in: in std_logic_vector(7 downto 0);
  user_senha: buffer std_logic_vector(7 downto 0);
  user_login: out std_logic_vector(3 downto 0);
  flag_senha, flag_admin: out std_logic
);
END Operativa;

ARCHITECTURE arq_Operativa OF Operativa IS
	
TYPE STATE_TYPE IS (HOLD, FUNC_SET, DISPLAY_ON, MODE_SET, WRITE_CHAR1,
WRITE_CHAR2,WRITE_CHAR3,WRITE_CHAR4,WRITE_CHAR5,WRITE_CHAR6,WRITE_CHAR7,
WRITE_CHAR8, WRITE_CHAR9, WRITE_CHAR10, WRITE_CHAR11, WRITE_CHAR12, 
WRITE_CHAR13, WRITE_CHAR14, WRITE_CHAR15, WRITE_CHAR16, RETURN_HOME, TOGGLE_E, RESET1, RESET2, 
RESET3, DISPLAY_OFF, DISPLAY_CLEAR);
SIGNAL state, next_command: STATE_TYPE;
SIGNAL DATA_BUS_VALUE: STD_LOGIC_VECTOR(7 DOWNTO 0);

SIGNAL CLK_COUNT_5HZ: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL CLK_5HZ : STD_LOGIC;
signal BCD_senha1, BCD_senha0: std_logic_vector(3 downto 0);
signal BCD_digit1, BCD_digit0, BCD_digit_aux: std_logic_vector(3 downto 0);

signal BCD_char1, BCD_char2, BCD_char3, BCD_char4, BCD_char5, BCD_char6, BCD_char7: std_logic_vector(7 downto 0);
signal BCD_char8, BCD_char9, BCD_char10, BCD_char11, BCD_char12, BCD_char13: std_logic_vector(7 downto 0);
signal BCD_char14, BCD_char15, BCD_char16: std_logic_vector(7 downto 0);
signal flag1_senha, flag2_admin: std_logic;
signal user_login1: std_logic_vector(3 downto 0);

BEGIN


  LCD_ON <= '1';
  RESET_LED <= not RESET;
  -- BIDIRECTIONAL TRI STATE LCD DATA BUS
  DATA_BUS <= DATA_BUS_VALUE WHEN LCD_RW = '0' ELSE "ZZZZZZZZ";


    
  PROCESS (clk, reset)
  BEGIN
    if reset = '0' then
	    state <= RESET1;
	    DATA_BUS_VALUE <= X"38";
	    next_command <= RESET2;
	    LCD_E <= '1';
	    LCD_RS <= '0';
	    LCD_RW <= '0';
	ELSIF clk'EVENT AND clk = '1' THEN
	
      IF CLK_COUNT_5HZ < 39 THEN
	    CLK_COUNT_5HZ <= CLK_COUNT_5HZ + 1;
	  ELSE
		CLK_COUNT_5HZ <= X"00";
		CLK_5HZ <= NOT CLK_5HZ;
	  END IF;

--casos LCD
	  CASE state IS
	    WHEN RESET1 =>
	      LCD_E <= '1';
		  LCD_RS <= '0';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= X"38";
		  state <= TOGGLE_E;
		  next_command <= RESET2;
		WHEN RESET2 =>
		  LCD_E <= '1';
		  LCD_RS <= '0';
		  LCD_RW <= '0';
	      DATA_BUS_VALUE <= X"38";
		  state <= TOGGLE_E;
		  next_command <= RESET3;
		WHEN RESET3 =>
		  LCD_E <= '1';
		  LCD_RS <= '0';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= X"38";
		  state <= TOGGLE_E;
		  next_command <= FUNC_SET;
-- EXTRA STATES ABOVE ARE NEEDED FOR RELIABLE PUSHBUTTON RESET OF LCD
		WHEN FUNC_SET =>
		  LCD_E <= '1';
		  LCD_RS <= '0';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= X"38";
		  state <= TOGGLE_E;
		  next_command <= DISPLAY_OFF;
-- Turn off Display and Turn off cursor
		WHEN DISPLAY_OFF =>
		  LCD_E <= '1';
		  LCD_RS <= '0';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= X"08";
		  state <= TOGGLE_E;
		  next_command <= DISPLAY_CLEAR;
-- Turn on Display and Turn off cursor
		WHEN DISPLAY_CLEAR =>
		  LCD_E <= '1';
		  LCD_RS <= '0';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= X"01";
		  state <= TOGGLE_E;
		  next_command <= DISPLAY_ON;
-- Turn on Display and Turn off cursor
		WHEN DISPLAY_ON =>
		  LCD_E <= '1';
		  LCD_RS <= '0';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= X"0C";
		  state <= TOGGLE_E;
		  next_command <= MODE_SET;
-- Set write mode to auto increment address and move cursor to the right
		WHEN MODE_SET =>
		  LCD_E <= '1';
		  LCD_RS <= '0';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= X"06";
		  state <= TOGGLE_E;
		  next_command <= WRITE_CHAR1;
-- Write ASCII hex character in first LCD character location
-- Um estado para cada caracter do LCD.
		WHEN WRITE_CHAR1 =>
		  LCD_E <= '1';
		  LCD_RS <= '1';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= BCD_char1;
		  state <= TOGGLE_E;
		  next_command <= WRITE_CHAR2;

		WHEN WRITE_CHAR2 =>
		  LCD_E <= '1';
		  LCD_RS <= '1';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= BCD_char2;
		  state <= TOGGLE_E;
		  next_command <= WRITE_CHAR3;

		WHEN WRITE_CHAR3 =>
		  LCD_E <= '1';
		  LCD_RS <= '1';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= BCD_char3;
		  state <= TOGGLE_E;
		  next_command <= WRITE_CHAR4;

		WHEN WRITE_CHAR4 =>
		  LCD_E <= '1';
		  LCD_RS <= '1';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= BCD_char4;
	      state <= TOGGLE_E;
		  next_command <= WRITE_CHAR5;

		WHEN WRITE_CHAR5 =>
		  LCD_E <= '1';
		  LCD_RS <= '1';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= BCD_char5;
		  state <= TOGGLE_E;
		  next_command <= WRITE_CHAR6;

		WHEN WRITE_CHAR6 =>
		  LCD_E <= '1';
		  LCD_RS <= '1';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= BCD_char6;
		  state <= TOGGLE_E;
		  next_command <= WRITE_CHAR7;

		WHEN WRITE_CHAR7 =>
		  LCD_E <= '1';
		  LCD_RS <= '1';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= BCD_char7;
		  state <= TOGGLE_E;
		  next_command <= WRITE_CHAR8;

		WHEN WRITE_CHAR8 =>
		  LCD_E <= '1';
		  LCD_RS <= '1';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= BCD_char8;
		  state <= TOGGLE_E;
		  next_command <= WRITE_CHAR9;

		WHEN WRITE_CHAR9 =>
		  LCD_E <= '1';
		  LCD_RS <= '1';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= BCD_char9;
		  state <= TOGGLE_E;
		  next_command <= WRITE_CHAR10;

		WHEN WRITE_CHAR10 =>
		  LCD_E <= '1';
		  LCD_RS <= '1';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= BCD_char10;
		  state <= TOGGLE_E;
		  next_command <= WRITE_CHAR11;

		WHEN WRITE_CHAR11 =>
		  LCD_E <= '1';
		  LCD_RS <= '1';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= BCD_char11;
		  state <= TOGGLE_E;
		  next_command <= WRITE_CHAR12;

		WHEN WRITE_CHAR12 =>
		  LCD_E <= '1';
		  LCD_RS <= '1';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= BCD_char12;
		  state <= TOGGLE_E;
		  next_command <= WRITE_CHAR13;

		WHEN WRITE_CHAR13 =>
		  LCD_E <= '1';
		  LCD_RS <= '1';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= BCD_char13;
		  state <= TOGGLE_E;
		  next_command <= WRITE_CHAR14;

		WHEN WRITE_CHAR14 =>
		  LCD_E <= '1';
		  LCD_RS <= '1';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= BCD_char14;
		  state <= TOGGLE_E;
		  next_command <= WRITE_CHAR15;

		WHEN WRITE_CHAR15 =>
		  LCD_E <= '1';
		  LCD_RS <= '1';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= BCD_char15;
		  state <= TOGGLE_E;
		  next_command <= WRITE_CHAR16;

		WHEN WRITE_CHAR16 =>
		  LCD_E <= '1';
		  LCD_RS <= '1';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= BCD_char16;
		  state <= TOGGLE_E;
		  next_command <= RETURN_HOME;

		WHEN RETURN_HOME =>
		  LCD_E <= '1';
		  LCD_RS <= '0';
		  LCD_RW <= '0';
		  DATA_BUS_VALUE <= X"80";
		  state <= TOGGLE_E;
	      next_command <= WRITE_CHAR1;
		
		WHEN TOGGLE_E =>
		  LCD_E <= '0';
		  state <= HOLD;

		WHEN HOLD =>
		  state <= next_command;
	  END CASE;
	END IF;
  END PROCESS;
  
--mensagens de cada estado no LCD.
  process(reset, clk)
  begin
    if reset='0' then
      BCD_char1 <= X"00";
      BCD_char2 <= X"00";
      BCD_char3 <= X"00";
      BCD_char4 <= X"00";
      BCD_char5 <= X"00";
      BCD_char6 <= X"00";
      BCD_char7 <= X"00";
      BCD_char8 <= X"00";
      BCD_char9 <= X"00";
      BCD_char10 <= X"00";
      BCD_char11 <= X"00";
      BCD_char12 <= X"00";
      BCD_char13 <= X"00";
      BCD_char14 <= X"00";
      BCD_char15 <= X"00";
      BCD_char16 <= X"00";
    elsif clk'event and clk='1' then
      if word_data_in="0000" then -- usuario;
		  BCD_char1 <= X"55";
		  BCD_char2 <= X"53";
		  BCD_char3 <= X"55";
		  BCD_char4 <= X"41";
		  BCD_char5 <= X"52";
		  BCD_char6 <= X"49";
		  BCD_char7 <= X"4F";
		  BCD_char8 <= X"3A";
		  BCD_char9 <= X"3" & BCD_digit1;
		  BCD_char10 <= X"3" & BCD_digit0;
		  BCD_char11 <= X"20";
		  BCD_char12 <= X"20";
		  BCD_char13 <= X"20";
		  BCD_char14 <= X"20";
		  BCD_char15 <= X"20";
		  BCD_char16 <= X"20"; 
      
      elsif word_data_in="0001" then -- senha;
		  BCD_char1 <= X"53";
		  BCD_char2 <= X"45";
		  BCD_char3 <= X"4E";
		  BCD_char4 <= X"48";
		  BCD_char5 <= X"41";
		  BCD_char6 <= X"3A";
		  BCD_char7 <= X"3" & BCD_senha1;
		  BCD_char8 <= X"3" & BCD_senha0;
		  BCD_char9 <= X"20";
		  BCD_char10 <= X"20";
		  BCD_char11 <= X"20";
		  BCD_char12 <= X"20";
		  BCD_char13 <= X"20";
		  BCD_char14 <= X"20";
		  BCD_char15 <= X"20";
		  BCD_char16 <= X"20";
		  
      elsif word_data_in="0010" then -- usuario invalido;
		  BCD_char1 <= X"55";
		  BCD_char2 <= X"53";
		  BCD_char3 <= X"55";
		  BCD_char4 <= X"41";
		  BCD_char5 <= X"52";
		  BCD_char6 <= X"49";
		  BCD_char7 <= X"4F";
		  BCD_char8 <= X"20";
		  BCD_char9 <= X"49";
		  BCD_char10 <= X"4E";
		  BCD_char11 <= X"56";
		  BCD_char12 <= X"41";
		  BCD_char13 <= X"4C";
		  BCD_char14 <= X"49";
		  BCD_char15 <= X"44";
		  BCD_char16 <= X"4F";
      
      elsif word_data_in="0011" then -- senha errada;
		  BCD_char1 <= X"53";
		  BCD_char2 <= X"45";
		  BCD_char3 <= X"4E";
		  BCD_char4 <= X"48";
		  BCD_char5 <= X"41";
		  BCD_char6 <= X"20";
		  BCD_char7 <= X"45";
		  BCD_char8 <= X"52";
		  BCD_char9 <= X"52";
		  BCD_char10 <= X"41";
		  BCD_char11 <= X"44";
		  BCD_char12 <= X"41";
		  BCD_char13 <= X"3A";
		  BCD_char14 <= X"20";
		  BCD_char15 <= X"20";
		  BCD_char16 <= X"20";
      
      elsif word_data_in="0100" then -- novo usuario;
		  BCD_char1 <= X"4E";
		  BCD_char2 <= X"4F";
		  BCD_char3 <= X"56";
		  BCD_char4 <= X"4F";
		  BCD_char5 <= X"20";
		  BCD_char6 <= X"55";
		  BCD_char7 <= X"53";
		  BCD_char8 <= X"55";
		  BCD_char9 <= X"41";
		  BCD_char10 <= X"52";
		  BCD_char11 <= X"49";
		  BCD_char12 <= X"4F";
		  BCD_char13 <= X"3A";
		  BCD_char14 <= X"3" & posicao1;
		  BCD_char15 <= X"3" & posicao0;
		  BCD_char16 <= X"20";
      
      elsif word_data_in="0101" then -- nova senha;
		  BCD_char1 <= X"4E";
		  BCD_char2 <= X"4F";
		  BCD_char3 <= X"56";
		  BCD_char4 <= X"41";
		  BCD_char5 <= X"20";
		  BCD_char6 <= X"53";
		  BCD_char7 <= X"45";
		  BCD_char8 <= X"4E";
		  BCD_char9 <= X"48";
		  BCD_char10 <= X"41";
		  BCD_char11 <= X"3A";
		  BCD_char12 <= X"3" & BCD_senha1;
		  BCD_char13 <= X"3" & BCD_senha0;
		  BCD_char14 <= X"20";
		  BCD_char15 <= X"20";
		  BCD_char16 <= X"20";
      
      elsif word_data_in="0110" then -- bem vindo;
		  BCD_char1 <= X"42";
		  BCD_char2 <= X"45";
		  BCD_char3 <= X"4D";
		  BCD_char4 <= X"20";
		  BCD_char5 <= X"56";
		  BCD_char6 <= X"49";
		  BCD_char7 <= X"4E";
		  BCD_char8 <= X"44";
		  BCD_char9 <= X"4F";
		  BCD_char10 <= X"20";
		  BCD_char11 <= X"20";
		  BCD_char12 <= X"20";
		  BCD_char13 <= X"20";
		  BCD_char14 <= X"20";
		  BCD_char15 <= X"20";
		  BCD_char16 <= X"20";
      
      else -- espere;
		  BCD_char1 <= X"45";
		  BCD_char2 <= X"53";
		  BCD_char3 <= X"50";
		  BCD_char4 <= X"45";
		  BCD_char5 <= X"52";
		  BCD_char6 <= X"45";
		  BCD_char7 <= X"20";
		  BCD_char8 <= X"20";
		  BCD_char9 <= X"20";
		  BCD_char10 <= X"20";
		  BCD_char11 <= X"20";
		  BCD_char12 <= X"20";
		  BCD_char13 <= X"20";
		  BCD_char14 <= X"20";
		  BCD_char15 <= X"20";
		  BCD_char16 <= X"20";
      end if;
    end if;
  end process;
  
--parte operativa senha.
  process(reset, CLK_5HZ)
  begin
    if reset='0' then
      BCD_senha1 <= X"0";
      BCD_senha0 <= X"0";
    elsif CLK_5HZ'event and CLK_5HZ='1' then
      if (btn1='0') then
        if BCD_senha1 < 9 then
          BCD_senha1 <= BCD_senha1 + 1;
        else
          BCD_senha1 <= X"0";
        end if;
      elsif (btn2='0') then
        if BCD_senha0 < 9 then
          BCD_senha0 <= BCD_senha0 + 1;
        else
          BCD_senha0 <= X"0";
        end if;
	  end if;
    end if;
    user_senha(3 downto 0) <= BCD_senha0;
    user_senha(7 downto 4) <= BCD_senha1;
  end process;
  
--parte operativa de login.
  process(reset, CLK_5HZ)
  begin
    if reset='0' then
      BCD_digit1 <= X"0";
      BCD_digit0 <= X"0";
      BCD_digit_aux <= X"0";
    elsif CLK_5HZ'event and CLK_5HZ='1' then
      if (btn2='0') then
	    BCD_digit0 <= BCD_digit0 + 1;
        BCD_digit_aux <= BCD_digit_aux + 1;
        if BCD_digit0=X"9" then
          BCD_digit0 <= X"0";
          BCD_digit1 <= BCD_digit1 + 1;
        elsif BCD_digit_aux=X"F" then
          BCD_digit0 <= X"0";
          BCD_digit1 <= X"0";
          BCD_digit_aux <= X"0";
        end if;
	  end if;
    end if;
    user_login1 <= BCD_digit_aux;
    user_login <= BCD_digit_aux;
  end process;
  
-- flags: login adm/user e senha.
  process(btn0)
  begin
    if btn0'event and btn0='0' then
      if user_login1=X"F" then
        flag2_admin <= '1';
      else
        flag2_admin <= '0';
      end if;
      
      if reg_data_in=user_senha then
        flag1_senha <= '1';
      else
        flag1_senha <= '0';
      end if;
    end if;
    flag_senha <= flag1_senha;
    flag_admin <= flag2_admin;
  end process;
  
END arq_Operativa;