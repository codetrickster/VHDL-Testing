LIBRARY	IEEE;
USE IEEE.std_logic_1164.all;

ENTITY seg15 IS
  PORT(
  ent: in std_logic_vector(7 downto 0);
  s: out std_logic_vector(20 downto 0)
  );
end seg15;
architecture arq_seg15 of seg15 is
begin 
  with ent select
  
  s <= "100000010000001000000" when "00000000",
       "100000010000001111001" when "00000001",
       "100000010000000100100" when "00000010",
       "100000010000000110000" when "00000011",
       "100000010000000011001" when "00000100",
       "100000010000000010010" when "00000101",
       "100000010000000000010" when "00000110",
       "100000010000001111000" when "00000111",
       "100000010000000000000" when "00001000",
       "100000010000000010000" when "00001001",
       
       "100000011110011000000" when "00001010",
       "100000011110011111001" when "00001011",
       "100000011110010100100" when "00001100",
       "100000011110010110000" when "00001101",
       "100000011110010011001" when "00001110",
       "100000011110010010010" when "00001111",
       "100000011110010000010" when "00010000",
       "100000011110011111000" when "00010001",
       "100000011110010000000" when "00010010",
       "100000011110010010000" when "00010011",
       
       "100000001001001000000" when "00010100",
       "100000001001001111001" when "00010101",
       "100000001001000100100" when "00010110",
       "100000001001000110000" when "00010111",
       "100000001001000011001" when "00011000",
       "100000001001000010010" when "00011001",
       "100000001001000000010" when "00011010",
       "100000001001001111000" when "00011011",
       "100000001001000000000" when "00011100",
       "100000001001000010000" when "00011101",
       
       "011111101111110111111" when others;
       
end arq_seg15;